magic
tech sky130A
timestamp 1733939897
<< nmos >>
rect -10 -25 5 25
<< ndiff >>
rect -45 15 -10 25
rect -45 -5 -40 15
rect -20 -5 -10 15
rect -45 -25 -10 -5
rect 5 15 40 25
rect 5 -5 15 15
rect 35 -5 40 15
rect 5 -25 40 -5
<< ndiffc >>
rect -40 -5 -20 15
rect 15 -5 35 15
<< psubdiff >>
rect -125 10 -75 25
rect -125 -10 -110 10
rect -90 -10 -75 10
rect -125 -25 -75 -10
<< psubdiffcont >>
rect -110 -10 -90 10
<< poly >>
rect -10 25 5 40
rect -10 -45 5 -25
rect -25 -50 20 -45
rect -25 -70 -15 -50
rect 10 -70 20 -50
rect -25 -75 20 -70
<< polycont >>
rect -15 -70 10 -50
<< locali >>
rect -125 15 -75 25
rect -45 15 -15 25
rect -125 10 -40 15
rect -125 -10 -110 10
rect -90 -5 -40 10
rect -20 -5 -15 15
rect -90 -10 -75 -5
rect -125 -25 -75 -10
rect -45 -25 -15 -5
rect 10 15 40 25
rect 10 -5 15 15
rect 35 -5 40 15
rect 10 -25 40 -5
rect -25 -50 20 -45
rect -25 -70 -15 -50
rect 10 -70 20 -50
rect -25 -75 20 -70
<< viali >>
rect -110 -10 -90 10
<< metal1 >>
rect -125 10 -75 25
rect -125 -10 -110 10
rect -90 -10 -75 10
rect -125 -25 -75 -10
<< labels >>
rlabel polycont -15 -70 10 -50 1 Input
rlabel poly -5 30 -5 30 1 Gate
rlabel metal1 -110 -10 -90 10 1 Ground
rlabel ndiffc -40 -5 -20 15 1 Source
rlabel ndiffc 15 -5 35 15 1 Drain
<< end >>
