* SPICE3 file created from pmos_sky130.ext - technology: sky130B

X0 Drain Input Vdd Vdd sky130_fd_pr__pfet_01v8 ad=0.2275 pd=2 as=0.2275 ps=2 w=0.65 l=0.15
